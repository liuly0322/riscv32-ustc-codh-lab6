
module mem #(                   //
        parameter  ADDR_LEN  = 11   //
    ) (
        input  clk, rst,
        input  [ADDR_LEN-1:0] addr, // memory address
        output reg [31:0] rd_data,  // data read out
        input  wr_req,
        input  [31:0] wr_data       // data write in
    );
    localparam MEM_SIZE = 1<<ADDR_LEN;
    reg [31:0] ram_cell [MEM_SIZE];

    always @ (posedge clk or posedge rst)
        if(rst)
            rd_data <= 0;
        else
            rd_data <= ram_cell[addr];

    always @ (posedge clk)
        if(wr_req)
            ram_cell[addr] <= wr_data;

endmodule
